magic
tech scmos
timestamp 1544200725
<< nwell >>
rect -24 -7 16 31
<< ntransistor >>
rect -13 -59 -11 -49
rect -5 -59 -3 -49
rect 3 -59 5 -49
<< ptransistor >>
rect -13 -1 -11 19
rect -5 -1 -3 19
rect 3 -1 5 19
<< ndiffusion >>
rect -14 -59 -13 -49
rect -11 -59 -10 -49
rect -6 -59 -5 -49
rect -3 -59 -2 -49
rect 2 -59 3 -49
rect 5 -59 6 -49
<< pdiffusion >>
rect -14 -1 -13 19
rect -11 -1 -10 19
rect -6 -1 -5 19
rect -3 -1 -2 19
rect 2 -1 3 19
rect 5 -1 6 19
<< ndcontact >>
rect -18 -59 -14 -49
rect -10 -59 -6 -49
rect -2 -59 2 -49
rect 6 -59 10 -49
<< pdcontact >>
rect -18 -1 -14 19
rect -10 -1 -6 19
rect -2 -1 2 19
rect 6 -1 10 19
<< psubstratepcontact >>
rect -18 -67 -14 -63
rect -6 -67 -2 -63
rect 6 -67 10 -63
<< nsubstratencontact >>
rect -18 23 -14 27
rect -6 23 -2 27
rect 6 23 10 27
<< polysilicon >>
rect -13 19 -11 21
rect -5 19 -3 21
rect 3 19 5 21
rect -13 -13 -11 -1
rect -13 -49 -11 -17
rect -5 -42 -3 -1
rect 3 -20 5 -1
rect -5 -49 -3 -46
rect 3 -49 5 -24
rect -13 -61 -11 -59
rect -5 -61 -3 -59
rect 3 -61 5 -59
<< polycontact >>
rect -15 -17 -11 -13
rect 1 -24 5 -20
rect -7 -46 -3 -42
<< metal1 >>
rect -21 27 13 28
rect -21 23 -18 27
rect -14 23 -6 27
rect -2 23 6 27
rect 10 23 13 27
rect -21 22 13 23
rect -18 19 -14 22
rect -2 19 2 22
rect -10 -6 -6 -1
rect 6 -13 10 -1
rect -18 -24 -10 -20
rect -6 -24 1 -20
rect -18 -49 -14 -24
rect 6 -49 10 -46
rect -2 -62 2 -59
rect -21 -63 13 -62
rect -21 -67 -18 -63
rect -14 -67 -6 -63
rect -2 -67 6 -63
rect 10 -67 13 -63
rect -21 -68 13 -67
<< m2contact >>
rect -10 -10 -6 -6
rect 6 -17 10 -13
rect -10 -24 -6 -20
rect 6 -46 10 -42
<< metal2 >>
rect -10 -20 -6 -10
rect 6 -42 10 -17
<< labels >>
rlabel polycontact -13 -15 -13 -15 3 A
rlabel metal1 -7 25 -7 25 5 vdd
rlabel polycontact -5 -44 -5 -44 1 B
rlabel metal1 -8 -65 -8 -65 1 gnd
rlabel metal1 8 -11 8 -11 1 Z
<< end >>
